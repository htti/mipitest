
`timescale 1ns/1ns
module	Mipi_Config
(
	input		[9:0]	LUT_INDEX,
	output	reg	[41:0]	LUT_DATA,
	output		[9:0]	LUT_SIZE
);

assign	LUT_SIZE = 10'd604;

//-----------------------------------------------------------------
/////////////////////	Config Data LUT	  //////////////////////////	
always@(*)
begin
	case(LUT_INDEX)
	//read
	0 :		LUT_DATA	=	{8'h0,2'b10,16'h0000, 16'h0};	//chip_version
	1 :		LUT_DATA	=	{8'h0,2'b10,16'h0001, 16'h0};	
	2 :		LUT_DATA	=	{8'h0,2'b10,16'h0002, 16'h0};   //revision_number
	3 :		LUT_DATA	=	{8'h0,2'b10,16'h0003, 16'h0};   //manufacture_id
	4 :		LUT_DATA	=	{8'h0,2'b10,16'h0004, 16'h0};   //smia_version
	//load otp read
	//delay 100
	
	//write 16bits reg
	
	5  : 		LUT_DATA	= 	{8'd100,2'b11,16'h301a, 16'h0019}; //reset register
	//delay 100
	6  : 		LUT_DATA	= 	{8'd100,2'b11,16'h301a, 16'h0218};
	//default 3R
	7  : 		LUT_DATA	= 	{8'h0,2'b11,16'h3042, 16'h0000};
	8  : 		LUT_DATA	= 	{8'h0,2'b11,16'h30c0, 16'h1810};
	9  : 		LUT_DATA	= 	{8'h0,2'b11,16'h30c8, 16'h0018};
	10 : 		LUT_DATA	= 	{8'h0,2'b11,16'h30d2, 16'h0000};
	11 : 		LUT_DATA	= 	{8'h0,2'b11,16'h30d4, 16'h3030};
	12 : 		LUT_DATA	= 	{8'h0,2'b11,16'h30d6, 16'h2200};
	13 : 		LUT_DATA	= 	{8'h0,2'b11,16'h30da, 16'h0080};
	14 : 		LUT_DATA	= 	{8'h0,2'b11,16'h30dc, 16'h0080};
	15 : 		LUT_DATA	= 	{8'h0,2'b11,16'h30ee, 16'h0340};
	16 : 		LUT_DATA	= 	{8'h0,2'b11,16'h316a, 16'h8800};
	17 : 		LUT_DATA	= 	{8'h0,2'b11,16'h316c, 16'h8200};
	18 : 		LUT_DATA	= 	{8'h0,2'b11,16'h316e, 16'h8200};
	19 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3172, 16'h0286};
	20 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3174, 16'h8000};
	21 : 		LUT_DATA	= 	{8'h0,2'b11,16'h317c, 16'hE103};
	22 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3180, 16'hB080};
	23 : 		LUT_DATA	= 	{8'h0,2'b11,16'h31e0, 16'h0741};
	24 : 		LUT_DATA	= 	{8'h0,2'b11,16'h31e6, 16'h0000};
	25 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3ecc, 16'h0056};
	26 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3ed0, 16'hA666};
	27 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3ed2, 16'h6664};
	28 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3ed4, 16'h6ACC};
	29 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3ed8, 16'h7488};
	30 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3eda, 16'h77CB};
	31 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3EDE, 16'h6664};
	32 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3EE0, 16'h26D5};
	
	33 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3EE4, 16'h3548};
	34 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3EE6, 16'hB10C};
	35 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3EE8, 16'h6E79};
	36 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3EEA, 16'hC8B9};
	37 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3EFA, 16'hA656};
	38 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3EFE, 16'h99CC};
	39 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F00, 16'h0028};
	40 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F02, 16'h0140};
	41 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F04, 16'h0002};
	42 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F06, 16'h0004};
	43 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F08, 16'h0008};
	44 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F0A, 16'h0B09};
	45 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F0C, 16'h0302};
	46 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F10, 16'h0505};
	47 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F12, 16'h0303};
	48 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F14, 16'h0101};
	49 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F16, 16'h2020};
	50 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F18, 16'h0404};
	51 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F1A, 16'h7070};
	52 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F1C, 16'h003A};
	53 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F1E, 16'h003C};
	54 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F20, 16'h0209};
	55 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F2C, 16'h2210};
	56 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F38, 16'h44A8};
	57 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F40, 16'h2020};
	58 : 		LUT_DATA	= 	{8'h0,2'b11,16'h3F42, 16'h0808};
	59 : 		LUT_DATA	= 	{8'd0,2'b11,16'h3F44, 16'h0101};
//	60 : 		LUT_DATA	= 	{8'h6c,2'b11,16'h3F18, 16'h26D5};
	//delay 100
	60  : 		LUT_DATA	= 	{8'd100,2'b10,16'h3D00, 16'h0400}; //HIGH 8BITS
	61  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D01, 16'h7100}; 
	62  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D02, 16'hC900}; 
	63  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D03, 16'hFF00}; 
	64  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D04, 16'hFF00}; 
	65  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D05, 16'hFF00}; 
	66  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D06, 16'hFF00}; 
	67  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D07, 16'hFF00}; 
	                                
	68  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D08, 16'h6F00}; 
	69  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D09, 16'h4000}; 
	70  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D0A, 16'h1400};
	71  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D0B, 16'h0E00};
	72  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D0C, 16'h2300};
	73  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D0D, 16'hC200};
	74  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D0E, 16'h4100};
	75  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D0F, 16'h2000};
	76  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D10, 16'h3000}; 
	77  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D11, 16'h5400}; 
	78  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D12, 16'h8000}; 
	79  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D13, 16'h4200};
	80  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D14, 16'h0000};
	81  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D15, 16'hC000};
	82  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D16, 16'h8300};
	83  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D17, 16'h5700};
	84  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D18, 16'h8400};
	85  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D19, 16'h6400};
	86  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D1A, 16'h6400};
	87  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D1B, 16'h5500};
	88  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D1C, 16'h8000};
	89  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D1D, 16'h2300};
	90  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D1E, 16'h0000};	
	91  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D1F, 16'h6500};
	92  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D20, 16'h6500};
	93  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D21, 16'h8200};
	94  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D22, 16'h0000};
	95  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D23, 16'hC000};
	96  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D24, 16'h6E00};
	97  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D25, 16'h8000};
	98  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D26, 16'h5000};
	99  : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D27, 16'h5100};
	100 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D28, 16'h8300};
	101 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D29, 16'h4200};
	102 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D2A, 16'h8300};
	103 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D2B, 16'h5800};
	104 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D2C, 16'h6E00};
	105 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D2D, 16'h8000};
	106 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D2E, 16'h5F00};	
	107 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D2F, 16'h8700};
	108 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D30, 16'h6300};
	109 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D31, 16'h8200};
	110 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D32, 16'h5B00};
	111 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D33, 16'h8200};
	112 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D34, 16'h5900};
	113 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D35, 16'h8000};
	114 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D36, 16'h5A00};
	115 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D37, 16'h5E00};
	116 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D38, 16'hBD00};
	117 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D39, 16'h5900};
	118 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D3A, 16'h5900};
	119 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D3B, 16'h9D00};
	120 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D3C, 16'h6C00};
	121 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D3D, 16'h8000};
	122 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D3E, 16'h6D00};
	123 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D3F, 16'hA300};
	124 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D40, 16'h5000};
	125 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D41, 16'h8000};
	126 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D42, 16'h5100};
	127 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D43, 16'h8200};
	128 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D44, 16'h5800};
	129 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D45, 16'h8000};
	130 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D46, 16'h6600};
	131 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D47, 16'h8300};
	132 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D48, 16'h6400};
	133 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D49, 16'h6400};
	134 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D4A, 16'h8000};
	135 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D4B, 16'h3000};
	136 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D4C, 16'h5000};
	137 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D4D, 16'hDC00};
	138 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D4E, 16'h6A00};
	139 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D4F, 16'h8300};
	140 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D50, 16'h6B00};
	141 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D51, 16'hAA00};
	142 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D52, 16'h3000};
	143 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D53, 16'h9400};
	144 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D54, 16'h6700};
	145 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D55, 16'h8400};
	146 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D56, 16'h6500};
	147 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D57, 16'h6500};
	148 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D58, 16'h8100};
	149 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D59, 16'h4D00};
	150 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D5A, 16'h6800};
	151 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D5B, 16'h6A00};
	152 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D5C, 16'hAC00};
	153 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D5D, 16'h0600};
	154 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D5E, 16'h0800};
	155 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D5F, 16'h8D00};
	156 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D60, 16'h4500};
	157 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D61, 16'h9600};
	158 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D62, 16'h4500};
	159 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D63, 16'h8500};
	160 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D64, 16'h6A00};
	161 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D65, 16'h8300};
	162 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D66, 16'h6B00};
	163 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D67, 16'h0600};
	164 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D68, 16'h0800};
	165 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D69, 16'hA900};
	166 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D6A, 16'h3000};
	167 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D6B, 16'h9000};
	168 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D6C, 16'h6700};
	169 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D6D, 16'h6400};
	170 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D6E, 16'h6400};
	171 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D6F, 16'h8900};
	172 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D70, 16'h6500};
	173 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D71, 16'h6500};
	174 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D72, 16'h8100};
	175 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D73, 16'h5800};
	176 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D74, 16'h8800};
	177 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D75, 16'h1000};
	178 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D76, 16'hC000};
	179 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D77, 16'hB100};
	180 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D78, 16'h5E00};
	181 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D79, 16'h9600};
	182 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D7A, 16'h5300};
	183 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D7B, 16'h8200};
	184 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D7C, 16'h5E00};
	185 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D7D, 16'h5200};
	186 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D7E, 16'h6600};
	187 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D7F, 16'h8000};
	188 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D80, 16'h5800};
	189 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D81, 16'h8300};
	190 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D82, 16'h6400};
	191 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D83, 16'h6400};
	192 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D84, 16'h8000};
	193 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D85, 16'h5B00};
	194 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D86, 16'h8100};
	195 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D87, 16'h5A00};
	196 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D88, 16'h1D00};
	197 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D89, 16'h0C00};
	198 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D8A, 16'h8000};
	199 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D8B, 16'h5500};
	200 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D8C, 16'h3000};
	201 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D8D, 16'h6000};
	202 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D8E, 16'h4100};
	203 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D8F, 16'h8200};
	204 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D90, 16'h4200};
	205 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D91, 16'hB200};
	206 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D92, 16'h4200};
	207 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D93, 16'h8000};
	208 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D94, 16'h4000};
	209 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D95, 16'h8100};
	210 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D96, 16'h4000};
	211 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D97, 16'h8900};
	212 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D98, 16'h0600};
	213 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D99, 16'hC000};
	214 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D9A, 16'h4100};
	215 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D9B, 16'h8000};
	216 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D9C, 16'h4200};
	217 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D9D, 16'h8500};
	218 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D9E, 16'h4400};
	219 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3D9F, 16'h8300};
	220 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA0, 16'h4300};
	221 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA1, 16'h8200};
	222 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA2, 16'h6A00};
	223 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA3, 16'h8300};
	224 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA4, 16'h6B00};
	225 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA5, 16'h8D00};
	226 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA6, 16'h4300};
	227 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA7, 16'h8300};
	228 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA8, 16'h4400};
	229 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DA9, 16'h8100};
	230 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DAA, 16'h4100};
	231 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DAB, 16'h8500};
	232 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DAC, 16'h0600};
	233 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DAD, 16'hC000};
	234 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DAE, 16'h8C00};
	235 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DAF, 16'h3000};
	236 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB0, 16'hA400};
	237 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB1, 16'h6700};
	238 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB2, 16'h8100};
	239 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB3, 16'h4200};
	240 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB4, 16'h8200};
	241 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB5, 16'h6500};
	242 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB6, 16'h6500};
	243 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB7, 16'h8100};
	244 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB8, 16'h6900};
	245 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DB9, 16'h6A00};
	246 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DBA, 16'h9600};
	247 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DBB, 16'h4000};
	248 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DBC, 16'h8200};
	249 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DBD, 16'h4000};
	250 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DBE, 16'h8900};
	251 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DBF, 16'h0600};
	252 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC0, 16'hC000};
	253 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC1, 16'h4100};
	254 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC2, 16'h8000};
	255 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC3, 16'h4200};
	256 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC4, 16'h8500};
	257 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC5, 16'h4400};
	258 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC6, 16'h8300};
	259 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC7, 16'h4300};
	260 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC8, 16'h9200};
	261 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DC9, 16'h4300};
	262 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DCA, 16'h8300};
	263 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DCB, 16'h4400};
	264 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DCC, 16'h8500};
	265 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DCD, 16'h4100};
	266 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DCE, 16'h8100};
	267 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DCF, 16'h0600};
	268 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD0, 16'hC000};
	269 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD1, 16'h8100};
	270 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD2, 16'h6A00};
	271 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD3, 16'h8300};
	272 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD4, 16'h6B00};
	273 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD5, 16'h8200};
	274 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD6, 16'h4200};
	275 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD7, 16'hA000};
	276 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD8, 16'h4000};
	277 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DD9, 16'h8400};
	278 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DDA, 16'h3800};
	279 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DDB, 16'hA800};
	280 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DDC, 16'h3300};
	281 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DDD, 16'h0000};
	282 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DDE, 16'h2800};
	283 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DDF, 16'h3000};
	284 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE0, 16'h7000};
	285 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE1, 16'h0000};
	286 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE2, 16'h6F00};
	287 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE3, 16'h4000};
	288 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE4, 16'h1400};
	289 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE5, 16'h0E00};
	290 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE6, 16'h2300};
	291 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE7, 16'hC200};
	292 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE8, 16'h4100};
	293 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DE9, 16'h8200};
	294 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DEA, 16'h4200};
	295 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DEB, 16'h0000};
	296 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DEC, 16'hC000};
	297 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DED, 16'h5D00};
	298 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DEE, 16'h8000};
	299 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DEF, 16'h5A00};
	300 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF0, 16'h8000};
	301 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF1, 16'h5700};
	302 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF2, 16'h8400};
	303 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF3, 16'h6400};
	304 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF4, 16'h8000};
	305 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF5, 16'h5500};
	306 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF6, 16'h8600};
	307 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF7, 16'h6400};
	308 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF8, 16'h8000};
	309 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DF9, 16'h6500};
	310 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DFA, 16'h8800};
	311 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DFB, 16'h6500};
	312 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DFC, 16'h8200};
	313 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DFD, 16'h5400};
	314 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DFE, 16'h8000};
	315 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3DFF, 16'h5800};
	316 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E00, 16'h8000};
	317 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E01, 16'h0000};
	318 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E02, 16'hC000};
	319 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E03, 16'h8600};
	320 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E04, 16'h4200};
	321 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E05, 16'h8200};
	322 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E06, 16'h1000};
	323 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E07, 16'h3000};
	324 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E08, 16'h9C00};
	325 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E09, 16'h5C00};
	326 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E0A, 16'h8000};
	327 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E0B, 16'h6E00};
	328 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E0C, 16'h8600};
	329 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E0D, 16'h5B00};
	330 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E0E, 16'h8000};
	331 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E0F, 16'h6300};
	332 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E10, 16'h9E00};
	333 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E11, 16'h5900};
	334 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E12, 16'h8C00};
	335 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E13, 16'h5E00};
	336 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E14, 16'h8A00};
	337 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E15, 16'h6C00};
	338 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E16, 16'h8000};
	339 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E17, 16'h6D00};
	340 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E18, 16'h8100};
	341 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E19, 16'h5F00};
	342 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E1A, 16'h6000};
	343 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E1B, 16'h6100};
	344 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E1C, 16'h8800};
	345 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E1D, 16'h1000};
	346 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E1E, 16'h3000};
	347 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E1F, 16'h6600};
	348 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E20, 16'h8300};
	349 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E21, 16'h6E00};
	350 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E22, 16'h8000};
	351 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E23, 16'h6400};
	352 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E24, 16'h8700};
	353 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E25, 16'h6400};
	354 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E26, 16'h3000};
	355 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E27, 16'h5000};
	356 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E28, 16'hD300};
	357 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E29, 16'h6A00};
	358 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E2A, 16'h6B00};
	359 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E2B, 16'hAD00};
	360 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E2C, 16'h3000};
	361 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E2D, 16'h9400};
	362 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E2E, 16'h6700};
	363 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E2F, 16'h8400};
	364 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E30, 16'h6500};
	365 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E31, 16'h8200};
	366 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E32, 16'h4D00};
	367 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E33, 16'h8300};
	368 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E34, 16'h6500};
	369 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E35, 16'h3000};
	370 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E36, 16'h5000};
	371 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E37, 16'hA700};
	372 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E38, 16'h4300};
	373 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E39, 16'h0600};
	374 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E3A, 16'h0000};
	375 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E3B, 16'h8D00};
	376 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E3C, 16'h4500};
	377 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E3D, 16'h9A00};
	378 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E3E, 16'h6A00};
	379 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E3F, 16'h6B00};
	380 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E40, 16'h4500};
	381 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E41, 16'h8500};
	382 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E42, 16'h0600};
	383 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E43, 16'h0000};
	384 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E44, 16'h8100};
	385 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E45, 16'h4300};
	386 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E46, 16'h8A00};
	387 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E47, 16'h6F00};
	388 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E48, 16'h9600};
	389 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E49, 16'h3000};
	390 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E4A, 16'h9000};
	391 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E4B, 16'h6700};
	392 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E4C, 16'h6400};
	393 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E4D, 16'h8800};
	394 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E4E, 16'h6400};
	395 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E4F, 16'h8000};
	396 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E50, 16'h6500};
	397 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E51, 16'h8200};
	398 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E52, 16'h1000};
	399 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E53, 16'hC000};
	400 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E54, 16'h8400};
	401 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E55, 16'h6500};
	402 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E56, 16'hEF00};
	403 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E57, 16'h1000};
	404 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E58, 16'hC000};
	405 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E59, 16'h6600};
	406 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E5A, 16'h8500};
	407 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E5B, 16'h6400};
	408 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E5C, 16'h8100};
	409 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E5D, 16'h1700};
	410 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E5E, 16'h0000};
	411 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E5F, 16'h8000};
	412 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E60, 16'h2000};
	413 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E61, 16'h0D00};
	414 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E62, 16'h8000};
	415 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E63, 16'h1800};
	416 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E64, 16'h0C00};
	417 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E65, 16'h8000};
	418 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E66, 16'h6400};
	419 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E67, 16'h3000};
	420 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E68, 16'h6000};
	421 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E69, 16'h4100};
	422 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E6A, 16'h8200};
	423 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E6B, 16'h4200};
	424 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E6C, 16'hB200};
	425 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E6D, 16'h4200};
	426 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E6E, 16'h8000};
	427 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E6F, 16'h4000};
	428 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E70, 16'h8200};
	429 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E71, 16'h4000};
	430 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E72, 16'h4C00};
	431 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E73, 16'h4500};
	432 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E74, 16'h9200};
	433 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E75, 16'h6A00};
	434 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E76, 16'h6B00};
	435 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E77, 16'h9B00};
	436 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E78, 16'h4500};
	437 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E79, 16'h8100};
	438 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E7A, 16'h4C00};
	439 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E7B, 16'h4000};
	440 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E7C, 16'h8C00};
	441 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E7D, 16'h3000};
	442 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E7E, 16'hA400};
	443 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E7F, 16'h6700};
	444 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E80, 16'h8500};
	445 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E81, 16'h6500};
	446 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E82, 16'h8700};
	447 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E83, 16'h6500};
	448 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E84, 16'h3000};
	449 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E85, 16'h6000};
	450 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E86, 16'hD300};
	451 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E87, 16'h6A00};
	452 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E88, 16'h6B00};
	453 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E89, 16'hAC00};
	454 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E8A, 16'h6C00};
	455 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E8B, 16'h3200};
	456 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E8C, 16'hA800};
	457 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E8D, 16'h8000};
	458 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E8E, 16'h2800};
	459 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E8F, 16'h3000};
	460 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E90, 16'h7000};
	461 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E91, 16'h0000};
	462 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E92, 16'h8000};
	463 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E93, 16'h4000};
	464 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E94, 16'h4C00};
	465 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E95, 16'hBD00};
	466 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E96, 16'h0000};
	467 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E97, 16'h0E00};
	468 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E98, 16'hBE00};
	469 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E99, 16'h4400};
	470 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E9A, 16'h8800};
	471 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E9B, 16'h4400};
	472 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E9C, 16'hBC00};
	473 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E9D, 16'h7800};
	474 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E9E, 16'h0900};
	475 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3E9F, 16'h0000};
	476 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA0, 16'h8900};
	477 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA1, 16'h0400};
	478 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA2, 16'h8000};
	479 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA3, 16'h8000};
	480 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA4, 16'h0200};
	481 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA5, 16'h4000};
	482 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA6, 16'h8600};
	483 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA7, 16'h0900};
	484 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA8, 16'h0000};
	485 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EA9, 16'h8E00};
	486 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EAA, 16'h0900};
	487 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EAB, 16'h0000};
	488 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EAC, 16'h8000};
	489 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EAD, 16'h0200};
	490 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EAE, 16'h4000};
	491 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EAF, 16'h8000};
	492 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB0, 16'h0400};
	493 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB1, 16'h8000};
	494 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB2, 16'h8800};
	495 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB3, 16'h7D00};
	496 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB4, 16'hA000};
	497 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB5, 16'h8600};
	498 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB6, 16'h0900};
	499 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB7, 16'h0000};
	500 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB8, 16'h8700};
	501 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EB9, 16'h7A00};
	502 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EBA, 16'h0000};
	503 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EBB, 16'h0E00};
	504 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EBC, 16'hC300};
	505 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EBD, 16'h7900};
	506 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EBE, 16'h4C00};
	507 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EBF, 16'h4000};
	508 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC0, 16'hBF00};
	509 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC1, 16'h7000};
	510 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC2, 16'h0000};
	511 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC3, 16'h0000};
	512 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC4, 16'h0000};
	513 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC5, 16'h0000};
	514 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC6, 16'h0000};
	515 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC7, 16'h0000};
	516 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC8, 16'h0000};
	517 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3EC9, 16'h0000};
	518 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3ECA, 16'h0000};
	519 : 		LUT_DATA	= 	{8'h0,2'b10,16'h3ECB, 16'h0000};	
	520	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0300, 16'h0005};          // VT_PIX_CLK_DIV
	521	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0302, 16'h0001};          // VT_SYS_CLK_DIV
	522	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0304, 16'h0004};          // PRE_PLL_CLK_DIV
	523	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0306, 16'h0046};          // PLL_MULTIPLIER
	524	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0308, 16'h000A};          // OP_PIX_CLK_DIV
	525	:		LUT_DATA 	= 	{8'h0,2'b11,16'h030A, 16'h0001};          // OP_SYS_CLK_DIV
	526	:		LUT_DATA 	= 	{8'd0,2'b11,16'h3064, 16'h7800};          // SMIA_TEST	
		//Delay = 1
	527	:		LUT_DATA 	= 	{8'd1,2'b11,16'h31B0, 16'h0060};          // FRAME_PREAMBLE 
	528	:		LUT_DATA 	= 	{8'h0,2'b11,16'h31B2, 16'h0042};          // LINE_PREAMBLE
	529	:		LUT_DATA 	= 	{8'h0,2'b11,16'h31B4, 16'h4C36};          // MIPI_TIMING_0
	530	:		LUT_DATA 	= 	{8'h0,2'b11,16'h31B6, 16'h5218};          // MIPI_TIMING_1
	531	:		LUT_DATA 	= 	{8'h0,2'b11,16'h31B8, 16'h404A};          // MIPI_TIMING_2
	532	:		LUT_DATA 	= 	{8'h0,2'b11,16'h31BA, 16'h028A};          // MIPI_TIMING_3
	533	:		LUT_DATA 	= 	{8'd0,2'b11,16'h31BC, 16'h0008};          // MIPI_TIMING_4	
		//Delay = 1
	534	:		LUT_DATA 	= 	{8'd1,2'b11,16'h0342, 16'h1000};          // LINE_LENGTH_PCK 
	535	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0340, 16'h0556};          // FRAME_LENGTH_LINES
	536	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0202, 16'h0500};          // COARSE_INTEGRATION_TIME
	537	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0344, 16'h0008};          // X_ADDR_START
	538	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0348, 16'h0CC5};          // X_ADDR_END
	539	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0346, 16'h0008};          // Y_ADDR_START
	540	:		LUT_DATA 	= 	{8'h0,2'b11,16'h034A, 16'h0995};          // Y_ADDR_END
	541	:		LUT_DATA 	= 	{8'h0,2'b11,16'h034C, 16'h0660};          // X_OUTPUT_SIZE
	542	:		LUT_DATA 	= 	{8'h0,2'b11,16'h034E, 16'h04C8};          // Y_OUTPUT_SIZE
	543	:		LUT_DATA 	= 	{8'h0,2'b11,16'h3040, 16'h68C3};          // READ_MODE
	544	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0400, 16'h0000};          // SCALING_MODE
	545	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0402, 16'h0000};          // SPATIAL_SAMPLING
	546	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0404, 16'h0010};          // SCALE_M
	547	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0408, 16'h1010};          // SECOND_RESIDUAL
	548	:		LUT_DATA 	= 	{8'h0,2'b11,16'h040A, 16'h0210};          // SECOND_CROP
	549	:		LUT_DATA 	= 	{8'h0,2'b11,16'h306E, 16'h9080};          // DATA_PATH_SELECT				
	550	:		LUT_DATA 	= 	{8'h0,2'b11,16'h301A, 16'h001C};          // RESET_REGISTER
		//[Go to Capture 3264 x 2448@15fps]
	551	:		LUT_DATA 	= 	{8'h0,2'b11,16'h301A, 16'h0218};          // RESET_REGISTER 				
	552	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0342, 16'h1000};     // LINE_LENGTH_PCK
	553	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0340, 16'h0AAC};    // FRAME_LENGTH_LINES
	554	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0202, 16'h0AAC};    // COARSE_INTEGRATION_TIME
	555	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0344, 16'h0008};     // X_ADDR_START
	556	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0348, 16'h0CC7};    // X_ADDR_END
	557	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0346, 16'h0008};     // Y_ADDR_START
	558	:		LUT_DATA 	= 	{8'h0,2'b11,16'h034A, 16'h0997};    // Y_ADDR_END
	559	:		LUT_DATA 	= 	{8'h0,2'b11,16'h034C, 16'h0CC0};    // X_OUTPUT_SIZE
	560	:		LUT_DATA 	= 	{8'h0,2'b11,16'h034E, 16'h0990};     // Y_OUTPUT_SIZE
	561	:		LUT_DATA 	= 	{8'h0,2'b11,16'h3040, 16'h4041};     // READ_MODE
	562	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0400, 16'h0000};     // SCALING_MODE
	563	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0402, 16'h0000};     // SPATIAL_SAMPLING
	564	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0404, 16'h0010};     // SCALE_M
	565	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0408, 16'h1010};     // SECOND_RESIDUAL
	566	:		LUT_DATA 	= 	{8'h0,2'b11,16'h040A, 16'h0210};    // SECOND_CROP
	567	:		LUT_DATA 	= 	{8'h0,2'b11,16'h306E, 16'h9080};     // DATA_PATH_SELECT
	568	:		LUT_DATA 	= 	{8'h0,2'b11,16'h301A, 16'h001C};    // RESET_REGISTER	
		//[Preview 1632 x 1224@30fps]
	569	:		LUT_DATA 	= 	{8'h0,2'b11,16'h301A, 16'h0218};          // RESET_REGISTER 				
	570	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0342, 16'h1000};          // LINE_LENGTH_PCK
	571	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0340, 16'h0556};          // FRAME_LENGTH_LINES
	572	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0202, 16'h0547};          // COARSE_INTEGRATION_TIME
	573	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0344, 16'h0008};          // X_ADDR_START
	574	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0348, 16'h0CC5};          // X_ADDR_END
	575	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0346, 16'h0008};          // Y_ADDR_START
	576	:		LUT_DATA 	= 	{8'h0,2'b11,16'h034A, 16'h0995};          // Y_ADDR_END
	577	:		LUT_DATA 	= 	{8'h0,2'b11,16'h034C, 16'h0660};          // X_OUTPUT_SIZE
	578	:		LUT_DATA 	= 	{8'h0,2'b11,16'h034E, 16'h04C8};          // Y_OUTPUT_SIZE
	579	:		LUT_DATA 	= 	{8'h0,2'b11,16'h3040, 16'h68C3};          // READ_MODE
	580	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0400, 16'h0000};          // SCALING_MODE
	581	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0402, 16'h0000};          // SPATIAL_SAMPLING
	582	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0404, 16'h0010};          // SCALE_M
	583	:		LUT_DATA 	= 	{8'h0,2'b11,16'h0408, 16'h1010};          // SECOND_RESIDUAL
	584	:		LUT_DATA 	= 	{8'h0,2'b11,16'h040A, 16'h0210};          // SECOND_CROP
	585	:		LUT_DATA 	= 	{8'h0,2'b11,16'h306E, 16'h9080};          // DATA_PATH_SELECT				
	586	:		LUT_DATA 	= 	{8'h0,2'b11,16'h301A, 16'h001C};          // RESET_REGISTER	
	                                                            
	587	:		LUT_DATA	= 	{8'h0,2'b10,16'h0101, 16'h0000};		//[Normal]								
	588	:		LUT_DATA	= 	{8'h0,2'b10,16'h0101, 16'h0100};       //[Horizontal Mirror]								
	589	:		LUT_DATA	= 	{8'h0,2'b10,16'h0101, 16'h0200};		//[Vertical Flip]								
	590	:		LUT_DATA	= 	{8'h0,2'b10,16'h0101, 16'h0300};		//[Rotate 180 degree]	
	                                                            
	591	:		LUT_DATA	= 	{8'h0,2'b11,16'h301A, 16'h0218}; // disable streaming [OTP read]
	592	:		LUT_DATA	= 	{8'h0,2'b11,16'h3134, 16'hCD95}; // timing parameters for otp read
	593	:		LUT_DATA	= 	{8'h0,2'b11,16'h3054, 16'h0400};				
	594	:		LUT_DATA	= 	{8'h0,2'b11,16'h304C, 16'h3000}; // choose to only read record type 0x30 //Record Type				
	595	:		LUT_DATA	= 	{8'h0,2'b11,16'h304A, 16'h0010}; // auto read start //Read Command
//read	                                                           
	596 :		LUT_DATA	=	{8'h10,2'b10,16'h0005,16'h0000};
	597 :		LUT_DATA	=	{8'h10,2'b10,16'h0006,16'h0000};
	598 :		LUT_DATA	=	{8'h10,2'b10,16'h0008,16'h0000};
	599 :		LUT_DATA	=	{8'h10,2'b10,16'h0009,16'h0000};
	600 :		LUT_DATA	=	{8'h10,2'b10,16'h3024,16'h0000};
	601 :		LUT_DATA	=	{8'h10,2'b10,16'h3025,16'h0000};
	602 :		LUT_DATA	=	{8'h10,2'b10,16'h0112,16'h0000};
	603 :		LUT_DATA	=	{8'h10,2'b10,16'h0113,16'h0000};
	
	default: LUT_DATA	=	{8'h0,2'b10,16'h1C, 16'h7F};
	endcase
	
end

endmodule
