`timescale 1ns/1ns
module	Mipi_Config1
(
	input		[9:0]	LUT_INDEX,
	output	reg	[41:0]	LUT_DATA,
	output		[9:0]	LUT_SIZE
);

assign	LUT_SIZE = 10'd583;

//-----------------------------------------------------------------
/////////////////////	Config Data LUT	  //////////////////////////	
always@(*)
begin
	case(LUT_INDEX)


//void BYD_CONFIG_1024x768_RAW8(bool bScale, bool bTestMode)
//{
//	printf("=====================================\r\n");
 //   printf("BYD_CONFIG, Scale=%s, TestMode=%s\r\n", bScale?"yes":"no", bTestMode?"yes":"no");
//	printf("=====================================\r\n");

    0   : LUT_DATA = { 8'd0  ,2'b11,16'h301A, 16'h0019}; 	// RESET_REGISTER
    1   : LUT_DATA = { 8'd100,2'b11,16'h301A, 16'h0218}; 	// RESET_REGISTER     Sleep(100);
    2   : LUT_DATA = { 8'd0  ,2'b11,16'h3042, 16'h0000}; 	// DARK_CONTROL2
    3   : LUT_DATA = { 8'd0  ,2'b11,16'h30C0, 16'h1810}; 	// CALIB_CONTROL
    4   : LUT_DATA = { 8'd0  ,2'b11,16'h30C8, 16'h0018}; 	// CALIB_DAC
    5   : LUT_DATA = { 8'd0  ,2'b11,16'h30D2, 16'h0000}; 	// CRM_CONTROL
    6   : LUT_DATA = { 8'd0  ,2'b11,16'h30D4, 16'hD030}; 	// COLUMN_CORRECTION
    7   : LUT_DATA = { 8'd0  ,2'b11,16'h30D6, 16'h2200}; 	// COLUMN_CORRECTION2
    8   : LUT_DATA = { 8'd0  ,2'b11,16'h30DA, 16'h0080}; 	// COLUMN_CORRECTION_CLIP2
    9   : LUT_DATA = { 8'd0  ,2'b11,16'h30DC, 16'h0080}; 	// COLUMN_CORRECTION_CLIP3
    10  : LUT_DATA = { 8'd0  ,2'b11,16'h30EE, 16'h0340}; 	// DARK_CONTROL3
    11  : LUT_DATA = { 8'd0  ,2'b11,16'h316A, 16'h8800}; 	// DAC_RSTLO
    12  : LUT_DATA = { 8'd0  ,2'b11,16'h316C, 16'h8200}; 	// DAC_TXLO
    13  : LUT_DATA = { 8'd0  ,2'b11,16'h3172, 16'h0286}; 	// ANALOG_CONTROL2
    14  : LUT_DATA = { 8'd0  ,2'b11,16'h3174, 16'h8000}; 	// ANALOG_CONTROL3
    15  : LUT_DATA = { 8'd0  ,2'b11,16'h317C, 16'hE103}; 	// ANALOG_CONTROL7
    16  : LUT_DATA = { 8'd0  ,2'b11,16'h3180, 16'hF0FF}; 	// FINEDIGCORR_CONTROL
    17  : LUT_DATA = { 8'd0  ,2'b11,16'h31E0, 16'h0741}; 	// PIX_DEF_ID
    18  : LUT_DATA = { 8'd0  ,2'b11,16'h3ECC, 16'h0056}; 	// DAC_LD_0_1
    19  : LUT_DATA = { 8'd0  ,2'b11,16'h3ED0, 16'hA8AA}; 	// DAC_LD_4_5
    20  : LUT_DATA = { 8'd0  ,2'b11,16'h3ED2, 16'hAAA8}; 	// DAC_LD_6_7
    21  : LUT_DATA = { 8'd0  ,2'b11,16'h3ED4, 16'h8ACC}; 	// DAC_LD_8_9
    22  : LUT_DATA = { 8'd0  ,2'b11,16'h3ED8, 16'h7288}; 	// DAC_LD_12_13
    23  : LUT_DATA = { 8'd0  ,2'b11,16'h3EDA, 16'h77CA}; 	// DAC_LD_14_15
    24  : LUT_DATA = { 8'd0  ,2'b11,16'h3EDE, 16'h6664}; 	// DAC_LD_18_19
    25  : LUT_DATA = { 8'd0  ,2'b11,16'h3EE0, 16'h26D5}; 	// DAC_LD_20_21
    26  : LUT_DATA = { 8'd0  ,2'b11,16'h3EE4, 16'h1548}; 	// DAC_LD_24_25
    27  : LUT_DATA = { 8'd0  ,2'b11,16'h3EE6, 16'hB10C}; 	// DAC_LD_26_27
    28  : LUT_DATA = { 8'd0  ,2'b11,16'h3EE8, 16'h6E79}; 	// DAC_LD_28_29
    29  : LUT_DATA = { 8'd0  ,2'b11,16'h3EFE, 16'h77CC}; 	// DAC_LD_TXLO
    30  : LUT_DATA = { 8'd0  ,2'b11,16'h31E6, 16'h0000}; 	// PIX_DEF_ID_2
    31  : LUT_DATA = { 8'd0  ,2'b11,16'h3F00, 16'h0028}; 	// BM_T0
    32  : LUT_DATA = { 8'd0  ,2'b11,16'h3F02, 16'h0140}; 	// BM_T1
    33  : LUT_DATA = { 8'd0  ,2'b11,16'h3F04, 16'h0002}; 	// NOISE_GAIN_THRESHOLD0
    34  : LUT_DATA = { 8'd0  ,2'b11,16'h3F06, 16'h0004}; 	// NOISE_GAIN_THRESHOLD1
    35  : LUT_DATA = { 8'd0  ,2'b11,16'h3F08, 16'h0008}; 	// NOISE_GAIN_THRESHOLD2
    36  : LUT_DATA = { 8'd0  ,2'b11,16'h3F0A, 16'h0B09}; 	// NOISE_FLOOR10
    37  : LUT_DATA = { 8'd0  ,2'b11,16'h3F0C, 16'h0302}; 	// NOISE_FLOOR32
    38  : LUT_DATA = { 8'd0  ,2'b11,16'h3F10, 16'h0505}; 	// SINGLE_K_FACTOR0
    39  : LUT_DATA = { 8'd0  ,2'b11,16'h3F12, 16'h0303}; 	// SINGLE_K_FACTOR1
    40  : LUT_DATA = { 8'd0  ,2'b11,16'h3F14, 16'h0101}; 	// SINGLE_K_FACTOR2
    41  : LUT_DATA = { 8'd0  ,2'b11,16'h3F16, 16'h2020}; 	// CROSSFACTOR0
    42  : LUT_DATA = { 8'd0  ,2'b11,16'h3F18, 16'h0404}; 	// CROSSFACTOR1
    43  : LUT_DATA = { 8'd0  ,2'b11,16'h3F1A, 16'h7070}; 	// CROSSFACTOR2
    44  : LUT_DATA = { 8'd0  ,2'b11,16'h3F1C, 16'h003A}; 	// SINGLE_MAXFACTOR
    45  : LUT_DATA = { 8'd0  ,2'b11,16'h3F1E, 16'h003C}; 	// NOISE_COEF
    46  : LUT_DATA = { 8'd0  ,2'b11,16'h3F2C, 16'h2210}; 	// GTH_THRES_RTN
    47  : LUT_DATA = { 8'd0  ,2'b11,16'h3F40, 16'h2020}; 	// COUPLE_K_FACTOR0
    48  : LUT_DATA = { 8'd0  ,2'b11,16'h3F42, 16'h0808}; 	// COUPLE_K_FACTOR1
    49  : LUT_DATA = { 8'd0  ,2'b11,16'h3F44, 16'h0101}; 	// COUPLE_K_FACTOR2
    50  : LUT_DATA = { 8'd100  ,2'b10,16'h3D00, 16'h0400};   //sleep 100
    51  : LUT_DATA = { 8'd0  ,2'b10,16'h3D01, 16'h7000};
    52  : LUT_DATA = { 8'd0  ,2'b10,16'h3D02, 16'hC800};
    53  : LUT_DATA = { 8'd0  ,2'b10,16'h3D03, 16'hFF00};
    54  : LUT_DATA = { 8'd0  ,2'b10,16'h3D04, 16'hFF00};
    55  : LUT_DATA = { 8'd0  ,2'b10,16'h3D05, 16'hFF00};
    56  : LUT_DATA = { 8'd0  ,2'b10,16'h3D06, 16'hFF00};
    57  : LUT_DATA = { 8'd0  ,2'b10,16'h3D07, 16'hFF00};
    58  : LUT_DATA = { 8'd0  ,2'b10,16'h3D08, 16'h6F00};
    59  : LUT_DATA = { 8'd0  ,2'b10,16'h3D09, 16'h4000};
    60  : LUT_DATA = { 8'd0  ,2'b10,16'h3D0A, 16'h1400};
    61  : LUT_DATA = { 8'd0  ,2'b10,16'h3D0B, 16'h0E00};
    62  : LUT_DATA = { 8'd0  ,2'b10,16'h3D0C, 16'h2300};
    63  : LUT_DATA = { 8'd0  ,2'b10,16'h3D0D, 16'h8200};
    64  : LUT_DATA = { 8'd0  ,2'b10,16'h3D0E, 16'h4100};
    65  : LUT_DATA = { 8'd0  ,2'b10,16'h3D0F, 16'h5C00};
    66  : LUT_DATA = { 8'd0  ,2'b10,16'h3D10, 16'h5400};
    67  : LUT_DATA = { 8'd0  ,2'b10,16'h3D11, 16'h6E00};
    68  : LUT_DATA = { 8'd0  ,2'b10,16'h3D12, 16'h4200};
    69  : LUT_DATA = { 8'd0  ,2'b10,16'h3D13, 16'h0000};
    70  : LUT_DATA = { 8'd0  ,2'b10,16'h3D14, 16'hC000};
    71  : LUT_DATA = { 8'd0  ,2'b10,16'h3D15, 16'h5D00};
    72  : LUT_DATA = { 8'd0  ,2'b10,16'h3D16, 16'h8000};
    73  : LUT_DATA = { 8'd0  ,2'b10,16'h3D17, 16'h5A00};
    74  : LUT_DATA = { 8'd0  ,2'b10,16'h3D18, 16'h8000};
    75  : LUT_DATA = { 8'd0  ,2'b10,16'h3D19, 16'h5700};
    76  : LUT_DATA = { 8'd0  ,2'b10,16'h3D1A, 16'h8400};
    77  : LUT_DATA = { 8'd0  ,2'b10,16'h3D1B, 16'h6400};
    78  : LUT_DATA = { 8'd0  ,2'b10,16'h3D1C, 16'h8000};
    79  : LUT_DATA = { 8'd0  ,2'b10,16'h3D1D, 16'h5500};
    80  : LUT_DATA = { 8'd0  ,2'b10,16'h3D1E, 16'h8600};
    81  : LUT_DATA = { 8'd0  ,2'b10,16'h3D1F, 16'h6400};
    82  : LUT_DATA = { 8'd0  ,2'b10,16'h3D20, 16'h8000};
    83  : LUT_DATA = { 8'd0  ,2'b10,16'h3D21, 16'h6500};
    84  : LUT_DATA = { 8'd0  ,2'b10,16'h3D22, 16'h8800};
    85  : LUT_DATA = { 8'd0  ,2'b10,16'h3D23, 16'h6500};
    86  : LUT_DATA = { 8'd0  ,2'b10,16'h3D24, 16'h8400};
    87  : LUT_DATA = { 8'd0  ,2'b10,16'h3D25, 16'h5800};
    88  : LUT_DATA = { 8'd0  ,2'b10,16'h3D26, 16'h8000};
    89  : LUT_DATA = { 8'd0  ,2'b10,16'h3D27, 16'h0000};
    90  : LUT_DATA = { 8'd0  ,2'b10,16'h3D28, 16'hC000};
    91  : LUT_DATA = { 8'd0  ,2'b10,16'h3D29, 16'h8000};
    92  : LUT_DATA = { 8'd0  ,2'b10,16'h3D2A, 16'h3000};
    93  : LUT_DATA = { 8'd0  ,2'b10,16'h3D2B, 16'h0C00};
    94  : LUT_DATA = { 8'd0  ,2'b10,16'h3D2C, 16'h8400};
    95  : LUT_DATA = { 8'd0  ,2'b10,16'h3D2D, 16'h4200};
    96  : LUT_DATA = { 8'd0  ,2'b10,16'h3D2E, 16'h8200};
    97  : LUT_DATA = { 8'd0  ,2'b10,16'h3D2F, 16'h1000};
    98  : LUT_DATA = { 8'd0  ,2'b10,16'h3D30, 16'h3000};
    99  : LUT_DATA = { 8'd0  ,2'b10,16'h3D31, 16'hA600};
    100 : LUT_DATA = { 8'd0  ,2'b10,16'h3D32, 16'h5B00};
    101 : LUT_DATA = { 8'd0  ,2'b10,16'h3D33, 16'h8000};
    102 : LUT_DATA = { 8'd0  ,2'b10,16'h3D34, 16'h6300};
    103 : LUT_DATA = { 8'd0  ,2'b10,16'h3D35, 16'h8B00};
    104 : LUT_DATA = { 8'd0  ,2'b10,16'h3D36, 16'h3000};
    105 : LUT_DATA = { 8'd0  ,2'b10,16'h3D37, 16'h0C00};
    106 : LUT_DATA = { 8'd0  ,2'b10,16'h3D38, 16'hA500};
    107 : LUT_DATA = { 8'd0  ,2'b10,16'h3D39, 16'h5900};
    108 : LUT_DATA = { 8'd0  ,2'b10,16'h3D3A, 16'h8400};
    109 : LUT_DATA = { 8'd0  ,2'b10,16'h3D3B, 16'h6C00};
    110 : LUT_DATA = { 8'd0  ,2'b10,16'h3D3C, 16'h8000};
    111 : LUT_DATA = { 8'd0  ,2'b10,16'h3D3D, 16'h6D00};
    112 : LUT_DATA = { 8'd0  ,2'b10,16'h3D3E, 16'h8100};
    113 : LUT_DATA = { 8'd0  ,2'b10,16'h3D3F, 16'h5F00};
    114 : LUT_DATA = { 8'd0  ,2'b10,16'h3D40, 16'h6000};
    115 : LUT_DATA = { 8'd0  ,2'b10,16'h3D41, 16'h6100};
    116 : LUT_DATA = { 8'd0  ,2'b10,16'h3D42, 16'h1000};
    117 : LUT_DATA = { 8'd0  ,2'b10,16'h3D43, 16'h3000};
    118 : LUT_DATA = { 8'd0  ,2'b10,16'h3D44, 16'h8800};
    119 : LUT_DATA = { 8'd0  ,2'b10,16'h3D45, 16'h6600};
    120 : LUT_DATA = { 8'd0  ,2'b10,16'h3D46, 16'h8300};
    121 : LUT_DATA = { 8'd0  ,2'b10,16'h3D47, 16'h6E00};
    122 : LUT_DATA = { 8'd0  ,2'b10,16'h3D48, 16'h8000};
    123 : LUT_DATA = { 8'd0  ,2'b10,16'h3D49, 16'h6400};
    124 : LUT_DATA = { 8'd0  ,2'b10,16'h3D4A, 16'h8700};
    125 : LUT_DATA = { 8'd0  ,2'b10,16'h3D4B, 16'h6400};
    126 : LUT_DATA = { 8'd0  ,2'b10,16'h3D4C, 16'h3000};
    127 : LUT_DATA = { 8'd0  ,2'b10,16'h3D4D, 16'h5000};
    128 : LUT_DATA = { 8'd0  ,2'b10,16'h3D4E, 16'hDA00};
    129 : LUT_DATA = { 8'd0  ,2'b10,16'h3D4F, 16'h6A00};
    130 : LUT_DATA = { 8'd0  ,2'b10,16'h3D50, 16'h8300};
    131 : LUT_DATA = { 8'd0  ,2'b10,16'h3D51, 16'h6B00};
    132 : LUT_DATA = { 8'd0  ,2'b10,16'h3D52, 16'hA600};
    133 : LUT_DATA = { 8'd0  ,2'b10,16'h3D53, 16'h3000};
    134 : LUT_DATA = { 8'd0  ,2'b10,16'h3D54, 16'h9400};
    135 : LUT_DATA = { 8'd0  ,2'b10,16'h3D55, 16'h6700};
    136 : LUT_DATA = { 8'd0  ,2'b10,16'h3D56, 16'h8400};
    137 : LUT_DATA = { 8'd0  ,2'b10,16'h3D57, 16'h6500};
    138 : LUT_DATA = { 8'd0  ,2'b10,16'h3D58, 16'h8200};
    139 : LUT_DATA = { 8'd0  ,2'b10,16'h3D59, 16'h4D00};
    140 : LUT_DATA = { 8'd0  ,2'b10,16'h3D5A, 16'h8300};
    141 : LUT_DATA = { 8'd0  ,2'b10,16'h3D5B, 16'h6500};
    142 : LUT_DATA = { 8'd0  ,2'b10,16'h3D5C, 16'h3000};
    143 : LUT_DATA = { 8'd0  ,2'b10,16'h3D5D, 16'h5000};
    144 : LUT_DATA = { 8'd0  ,2'b10,16'h3D5E, 16'hA600};
    145 : LUT_DATA = { 8'd0  ,2'b10,16'h3D5F, 16'h5800};
    146 : LUT_DATA = { 8'd0  ,2'b10,16'h3D60, 16'h4300};
    147 : LUT_DATA = { 8'd0  ,2'b10,16'h3D61, 16'h0600};
    148 : LUT_DATA = { 8'd0  ,2'b10,16'h3D62, 16'h0000};
    149 : LUT_DATA = { 8'd0  ,2'b10,16'h3D63, 16'h8D00};
    150 : LUT_DATA = { 8'd0  ,2'b10,16'h3D64, 16'h4500};
    151 : LUT_DATA = { 8'd0  ,2'b10,16'h3D65, 16'hA000};
    152 : LUT_DATA = { 8'd0  ,2'b10,16'h3D66, 16'h4500};
    153 : LUT_DATA = { 8'd0  ,2'b10,16'h3D67, 16'h6A00};
    154 : LUT_DATA = { 8'd0  ,2'b10,16'h3D68, 16'h8300};
    155 : LUT_DATA = { 8'd0  ,2'b10,16'h3D69, 16'h6B00};
    156 : LUT_DATA = { 8'd0  ,2'b10,16'h3D6A, 16'h0600};
    157 : LUT_DATA = { 8'd0  ,2'b10,16'h3D6B, 16'h0000};
    158 : LUT_DATA = { 8'd0  ,2'b10,16'h3D6C, 16'h8100};
    159 : LUT_DATA = { 8'd0  ,2'b10,16'h3D6D, 16'h4300};
    160 : LUT_DATA = { 8'd0  ,2'b10,16'h3D6E, 16'h9C00};
    161 : LUT_DATA = { 8'd0  ,2'b10,16'h3D6F, 16'h5800};
    162 : LUT_DATA = { 8'd0  ,2'b10,16'h3D70, 16'h8400};
    163 : LUT_DATA = { 8'd0  ,2'b10,16'h3D71, 16'h3000};
    164 : LUT_DATA = { 8'd0  ,2'b10,16'h3D72, 16'h9000};
    165 : LUT_DATA = { 8'd0  ,2'b10,16'h3D73, 16'h6700};
    166 : LUT_DATA = { 8'd0  ,2'b10,16'h3D74, 16'h6400};
    167 : LUT_DATA = { 8'd0  ,2'b10,16'h3D75, 16'h8800};
    168 : LUT_DATA = { 8'd0  ,2'b10,16'h3D76, 16'h6400};
    169 : LUT_DATA = { 8'd0  ,2'b10,16'h3D77, 16'h8000};
    170 : LUT_DATA = { 8'd0  ,2'b10,16'h3D78, 16'h6500};
    171 : LUT_DATA = { 8'd0  ,2'b10,16'h3D79, 16'h8800};
    172 : LUT_DATA = { 8'd0  ,2'b10,16'h3D7A, 16'h6500};
    173 : LUT_DATA = { 8'd0  ,2'b10,16'h3D7B, 16'h8200};
    174 : LUT_DATA = { 8'd0  ,2'b10,16'h3D7C, 16'h1000};
    175 : LUT_DATA = { 8'd0  ,2'b10,16'h3D7D, 16'hC000};
    176 : LUT_DATA = { 8'd0  ,2'b10,16'h3D7E, 16'hEB00};
    177 : LUT_DATA = { 8'd0  ,2'b10,16'h3D7F, 16'h1000};
    178 : LUT_DATA = { 8'd0  ,2'b10,16'h3D80, 16'hC000};
    179 : LUT_DATA = { 8'd0  ,2'b10,16'h3D81, 16'h6600};
    180 : LUT_DATA = { 8'd0  ,2'b10,16'h3D82, 16'h8500};
    181 : LUT_DATA = { 8'd0  ,2'b10,16'h3D83, 16'h6400};
    182 : LUT_DATA = { 8'd0  ,2'b10,16'h3D84, 16'h8100};
    183 : LUT_DATA = { 8'd0  ,2'b10,16'h3D85, 16'h1700};
    184 : LUT_DATA = { 8'd0  ,2'b10,16'h3D86, 16'h0000};
    185 : LUT_DATA = { 8'd0  ,2'b10,16'h3D87, 16'h8000};
    186 : LUT_DATA = { 8'd0  ,2'b10,16'h3D88, 16'h2000};
    187 : LUT_DATA = { 8'd0  ,2'b10,16'h3D89, 16'h0D00};
    188 : LUT_DATA = { 8'd0  ,2'b10,16'h3D8A, 16'h8000};
    189 : LUT_DATA = { 8'd0  ,2'b10,16'h3D8B, 16'h1800};
    190 : LUT_DATA = { 8'd0  ,2'b10,16'h3D8C, 16'h0C00};
    191 : LUT_DATA = { 8'd0  ,2'b10,16'h3D8D, 16'h8000};
    192 : LUT_DATA = { 8'd0  ,2'b10,16'h3D8E, 16'h6400};
    193 : LUT_DATA = { 8'd0  ,2'b10,16'h3D8F, 16'h3000};
    194 : LUT_DATA = { 8'd0  ,2'b10,16'h3D90, 16'h6000};
    195 : LUT_DATA = { 8'd0  ,2'b10,16'h3D91, 16'h4100};
    196 : LUT_DATA = { 8'd0  ,2'b10,16'h3D92, 16'h8200};
    197 : LUT_DATA = { 8'd0  ,2'b10,16'h3D93, 16'h4200};
    198 : LUT_DATA = { 8'd0  ,2'b10,16'h3D94, 16'hB200};
    199 : LUT_DATA = { 8'd0  ,2'b10,16'h3D95, 16'h4200};
    200 : LUT_DATA = { 8'd0  ,2'b10,16'h3D96, 16'h8000};
    201 : LUT_DATA = { 8'd0  ,2'b10,16'h3D97, 16'h4000};
    202 : LUT_DATA = { 8'd0  ,2'b10,16'h3D98, 16'h8100};
    203 : LUT_DATA = { 8'd0  ,2'b10,16'h3D99, 16'h4000};
    204 : LUT_DATA = { 8'd0  ,2'b10,16'h3D9A, 16'h8000};
    205 : LUT_DATA = { 8'd0  ,2'b10,16'h3D9B, 16'h4100};
    206 : LUT_DATA = { 8'd0  ,2'b10,16'h3D9C, 16'h8000};
    207 : LUT_DATA = { 8'd0  ,2'b10,16'h3D9D, 16'h4200};
    208 : LUT_DATA = { 8'd0  ,2'b10,16'h3D9E, 16'h8000};
    209 : LUT_DATA = { 8'd0  ,2'b10,16'h3D9F, 16'h4300};
    210 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA0, 16'h8300};
    211 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA1, 16'h0600};
    212 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA2, 16'hC000};
    213 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA3, 16'h8800};
    214 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA4, 16'h4400};
    215 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA5, 16'h8700};
    216 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA6, 16'h6A00};
    217 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA7, 16'h8300};
    218 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA8, 16'h6B00};
    219 : LUT_DATA = { 8'd0  ,2'b10,16'h3DA9, 16'h9200};
    220 : LUT_DATA = { 8'd0  ,2'b10,16'h3DAA, 16'h4400};
    221 : LUT_DATA = { 8'd0  ,2'b10,16'h3DAB, 16'h8800};
    222 : LUT_DATA = { 8'd0  ,2'b10,16'h3DAC, 16'h0600};
    223 : LUT_DATA = { 8'd0  ,2'b10,16'h3DAD, 16'hC800};
    224 : LUT_DATA = { 8'd0  ,2'b10,16'h3DAE, 16'h8100};
    225 : LUT_DATA = { 8'd0  ,2'b10,16'h3DAF, 16'h4100};
    226 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB0, 16'h8500};
    227 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB1, 16'h3000};
    228 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB2, 16'hA400};
    229 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB3, 16'h6700};
    230 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB4, 16'h8500};
    231 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB5, 16'h6500};
    232 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB6, 16'h8700};
    233 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB7, 16'h6500};
    234 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB8, 16'h3000};
    235 : LUT_DATA = { 8'd0  ,2'b10,16'h3DB9, 16'h6000};
    236 : LUT_DATA = { 8'd0  ,2'b10,16'h3DBA, 16'h8D00};
    237 : LUT_DATA = { 8'd0  ,2'b10,16'h3DBB, 16'h4200};
    238 : LUT_DATA = { 8'd0  ,2'b10,16'h3DBC, 16'h8200};
    239 : LUT_DATA = { 8'd0  ,2'b10,16'h3DBD, 16'h4000};
    240 : LUT_DATA = { 8'd0  ,2'b10,16'h3DBE, 16'h8200};
    241 : LUT_DATA = { 8'd0  ,2'b10,16'h3DBF, 16'h4000};
    242 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC0, 16'h8000};
    243 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC1, 16'h4100};
    244 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC2, 16'h8000};
    245 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC3, 16'h4200};
    246 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC4, 16'h8000};
    247 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC5, 16'h4300};
    248 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC6, 16'h8300};
    249 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC7, 16'h0600};
    250 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC8, 16'hC000};
    251 : LUT_DATA = { 8'd0  ,2'b10,16'h3DC9, 16'h8800};
    252 : LUT_DATA = { 8'd0  ,2'b10,16'h3DCA, 16'h4400};
    253 : LUT_DATA = { 8'd0  ,2'b10,16'h3DCB, 16'h9C00};
    254 : LUT_DATA = { 8'd0  ,2'b10,16'h3DCC, 16'h4400};
    255 : LUT_DATA = { 8'd0  ,2'b10,16'h3DCD, 16'h8800};
    256 : LUT_DATA = { 8'd0  ,2'b10,16'h3DCE, 16'h0600};
    257 : LUT_DATA = { 8'd0  ,2'b10,16'h3DCF, 16'hC800};
    258 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD0, 16'h8500};
    259 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD1, 16'h4100};
    260 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD2, 16'h6A00};
    261 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD3, 16'h8300};
    262 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD4, 16'h6B00};
    263 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD5, 16'hA000};
    264 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD6, 16'h4200};
    265 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD7, 16'h8200};
    266 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD8, 16'h4000};
    267 : LUT_DATA = { 8'd0  ,2'b10,16'h3DD9, 16'h6C00};
    268 : LUT_DATA = { 8'd0  ,2'b10,16'h3DDA, 16'h3A00};
    269 : LUT_DATA = { 8'd0  ,2'b10,16'h3DDB, 16'hA800};
    270 : LUT_DATA = { 8'd0  ,2'b10,16'h3DDC, 16'h8000};
    271 : LUT_DATA = { 8'd0  ,2'b10,16'h3DDD, 16'h2800};
    272 : LUT_DATA = { 8'd0  ,2'b10,16'h3DDE, 16'h3000};
    273 : LUT_DATA = { 8'd0  ,2'b10,16'h3DDF, 16'h7000};
    274 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE0, 16'h6F00};
    275 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE1, 16'h4000};
    276 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE2, 16'h1400};
    277 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE3, 16'h0E00};
    278 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE4, 16'h2300};
    279 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE5, 16'hC200};
    280 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE6, 16'h4100};
    281 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE7, 16'h8200};
    282 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE8, 16'h4200};
    283 : LUT_DATA = { 8'd0  ,2'b10,16'h3DE9, 16'h0000};
    284 : LUT_DATA = { 8'd0  ,2'b10,16'h3DEA, 16'hC000};
    285 : LUT_DATA = { 8'd0  ,2'b10,16'h3DEB, 16'h5D00};
    286 : LUT_DATA = { 8'd0  ,2'b10,16'h3DEC, 16'h8000};
    287 : LUT_DATA = { 8'd0  ,2'b10,16'h3DED, 16'h5A00};
    288 : LUT_DATA = { 8'd0  ,2'b10,16'h3DEE, 16'h8000};
    289 : LUT_DATA = { 8'd0  ,2'b10,16'h3DEF, 16'h5700};
    290 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF0, 16'h8400};
    291 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF1, 16'h6400};
    292 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF2, 16'h8000};
    293 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF3, 16'h5500};
    294 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF4, 16'h8600};
    295 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF5, 16'h6400};
    296 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF6, 16'h8000};
    297 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF7, 16'h6500};
    298 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF8, 16'h8800};
    299 : LUT_DATA = { 8'd0  ,2'b10,16'h3DF9, 16'h6500};
    300 : LUT_DATA = { 8'd0  ,2'b10,16'h3DFA, 16'h8200};
    301 : LUT_DATA = { 8'd0  ,2'b10,16'h3DFB, 16'h5400};
    302 : LUT_DATA = { 8'd0  ,2'b10,16'h3DFC, 16'h8000};
    303 : LUT_DATA = { 8'd0  ,2'b10,16'h3DFD, 16'h5800};
    304 : LUT_DATA = { 8'd0  ,2'b10,16'h3DFE, 16'h8000};
    305 : LUT_DATA = { 8'd0  ,2'b10,16'h3DFF, 16'h0000};
    306 : LUT_DATA = { 8'd0  ,2'b10,16'h3E00, 16'hC000};
    307 : LUT_DATA = { 8'd0  ,2'b10,16'h3E01, 16'h8600};
    308 : LUT_DATA = { 8'd0  ,2'b10,16'h3E02, 16'h4200};
    309 : LUT_DATA = { 8'd0  ,2'b10,16'h3E03, 16'h8200};
    310 : LUT_DATA = { 8'd0  ,2'b10,16'h3E04, 16'h1000};
    311 : LUT_DATA = { 8'd0  ,2'b10,16'h3E05, 16'h3000};
    312 : LUT_DATA = { 8'd0  ,2'b10,16'h3E06, 16'h9C00};
    313 : LUT_DATA = { 8'd0  ,2'b10,16'h3E07, 16'h5C00};
    314 : LUT_DATA = { 8'd0  ,2'b10,16'h3E08, 16'h8000};
    315 : LUT_DATA = { 8'd0  ,2'b10,16'h3E09, 16'h6E00};
    316 : LUT_DATA = { 8'd0  ,2'b10,16'h3E0A, 16'h8600};
    317 : LUT_DATA = { 8'd0  ,2'b10,16'h3E0B, 16'h5B00};
    318 : LUT_DATA = { 8'd0  ,2'b10,16'h3E0C, 16'h8000};
    319 : LUT_DATA = { 8'd0  ,2'b10,16'h3E0D, 16'h6300};
    320 : LUT_DATA = { 8'd0  ,2'b10,16'h3E0E, 16'h9E00};
    321 : LUT_DATA = { 8'd0  ,2'b10,16'h3E0F, 16'h5900};
    322 : LUT_DATA = { 8'd0  ,2'b10,16'h3E10, 16'h8C00};
    323 : LUT_DATA = { 8'd0  ,2'b10,16'h3E11, 16'h5E00};
    324 : LUT_DATA = { 8'd0  ,2'b10,16'h3E12, 16'h8A00};
    325 : LUT_DATA = { 8'd0  ,2'b10,16'h3E13, 16'h6C00};
    326 : LUT_DATA = { 8'd0  ,2'b10,16'h3E14, 16'h8000};
    327 : LUT_DATA = { 8'd0  ,2'b10,16'h3E15, 16'h6D00};
    328 : LUT_DATA = { 8'd0  ,2'b10,16'h3E16, 16'h8100};
    329 : LUT_DATA = { 8'd0  ,2'b10,16'h3E17, 16'h5F00};
    330 : LUT_DATA = { 8'd0  ,2'b10,16'h3E18, 16'h6000};
    331 : LUT_DATA = { 8'd0  ,2'b10,16'h3E19, 16'h6100};
    332 : LUT_DATA = { 8'd0  ,2'b10,16'h3E1A, 16'h8800};
    333 : LUT_DATA = { 8'd0  ,2'b10,16'h3E1B, 16'h1000};
    334 : LUT_DATA = { 8'd0  ,2'b10,16'h3E1C, 16'h3000};
    335 : LUT_DATA = { 8'd0  ,2'b10,16'h3E1D, 16'h6600};
    336 : LUT_DATA = { 8'd0  ,2'b10,16'h3E1E, 16'h8300};
    337 : LUT_DATA = { 8'd0  ,2'b10,16'h3E1F, 16'h6E00};
    338 : LUT_DATA = { 8'd0  ,2'b10,16'h3E20, 16'h8000};
    339 : LUT_DATA = { 8'd0  ,2'b10,16'h3E21, 16'h6400};
    340 : LUT_DATA = { 8'd0  ,2'b10,16'h3E22, 16'h8700};
    341 : LUT_DATA = { 8'd0  ,2'b10,16'h3E23, 16'h6400};
    342 : LUT_DATA = { 8'd0  ,2'b10,16'h3E24, 16'h3000};
    343 : LUT_DATA = { 8'd0  ,2'b10,16'h3E25, 16'h5000};
    344 : LUT_DATA = { 8'd0  ,2'b10,16'h3E26, 16'hD300};
    345 : LUT_DATA = { 8'd0  ,2'b10,16'h3E27, 16'h6A00};
    346 : LUT_DATA = { 8'd0  ,2'b10,16'h3E28, 16'h6B00};
    347 : LUT_DATA = { 8'd0  ,2'b10,16'h3E29, 16'hAD00};
    348 : LUT_DATA = { 8'd0  ,2'b10,16'h3E2A, 16'h3000};
    349 : LUT_DATA = { 8'd0  ,2'b10,16'h3E2B, 16'h9400};
    350 : LUT_DATA = { 8'd0  ,2'b10,16'h3E2C, 16'h6700};
    351 : LUT_DATA = { 8'd0  ,2'b10,16'h3E2D, 16'h8400};
    352 : LUT_DATA = { 8'd0  ,2'b10,16'h3E2E, 16'h6500};
    353 : LUT_DATA = { 8'd0  ,2'b10,16'h3E2F, 16'h8200};
    354 : LUT_DATA = { 8'd0  ,2'b10,16'h3E30, 16'h4D00};
    355 : LUT_DATA = { 8'd0  ,2'b10,16'h3E31, 16'h8300};
    356 : LUT_DATA = { 8'd0  ,2'b10,16'h3E32, 16'h6500};
    357 : LUT_DATA = { 8'd0  ,2'b10,16'h3E33, 16'h3000};
    358 : LUT_DATA = { 8'd0  ,2'b10,16'h3E34, 16'h5000};
    359 : LUT_DATA = { 8'd0  ,2'b10,16'h3E35, 16'hA700};
    360 : LUT_DATA = { 8'd0  ,2'b10,16'h3E36, 16'h4300};
    361 : LUT_DATA = { 8'd0  ,2'b10,16'h3E37, 16'h0600};
    362 : LUT_DATA = { 8'd0  ,2'b10,16'h3E38, 16'h0000};
    363 : LUT_DATA = { 8'd0  ,2'b10,16'h3E39, 16'h8D00};
    364 : LUT_DATA = { 8'd0  ,2'b10,16'h3E3A, 16'h4500};
    365 : LUT_DATA = { 8'd0  ,2'b10,16'h3E3B, 16'h9A00};
    366 : LUT_DATA = { 8'd0  ,2'b10,16'h3E3C, 16'h6A00};
    367 : LUT_DATA = { 8'd0  ,2'b10,16'h3E3D, 16'h6B00};
    368 : LUT_DATA = { 8'd0  ,2'b10,16'h3E3E, 16'h4500};
    369 : LUT_DATA = { 8'd0  ,2'b10,16'h3E3F, 16'h8500};
    370 : LUT_DATA = { 8'd0  ,2'b10,16'h3E40, 16'h0600};
    371 : LUT_DATA = { 8'd0  ,2'b10,16'h3E41, 16'h0000};
    372 : LUT_DATA = { 8'd0  ,2'b10,16'h3E42, 16'h8100};
    373 : LUT_DATA = { 8'd0  ,2'b10,16'h3E43, 16'h4300};
    374 : LUT_DATA = { 8'd0  ,2'b10,16'h3E44, 16'h8A00};
    375 : LUT_DATA = { 8'd0  ,2'b10,16'h3E45, 16'h6F00};
    376 : LUT_DATA = { 8'd0  ,2'b10,16'h3E46, 16'h9600};
    377 : LUT_DATA = { 8'd0  ,2'b10,16'h3E47, 16'h3000};
    378 : LUT_DATA = { 8'd0  ,2'b10,16'h3E48, 16'h9000};
    379 : LUT_DATA = { 8'd0  ,2'b10,16'h3E49, 16'h6700};
    380 : LUT_DATA = { 8'd0  ,2'b10,16'h3E4A, 16'h6400};
    381 : LUT_DATA = { 8'd0  ,2'b10,16'h3E4B, 16'h8800};
    382 : LUT_DATA = { 8'd0  ,2'b10,16'h3E4C, 16'h6400};
    383 : LUT_DATA = { 8'd0  ,2'b10,16'h3E4D, 16'h8000};
    384 : LUT_DATA = { 8'd0  ,2'b10,16'h3E4E, 16'h6500};
    385 : LUT_DATA = { 8'd0  ,2'b10,16'h3E4F, 16'h8200};
    386 : LUT_DATA = { 8'd0  ,2'b10,16'h3E50, 16'h1000};
    387 : LUT_DATA = { 8'd0  ,2'b10,16'h3E51, 16'hC000};
    388 : LUT_DATA = { 8'd0  ,2'b10,16'h3E52, 16'h8400};
    389 : LUT_DATA = { 8'd0  ,2'b10,16'h3E53, 16'h6500};
    390 : LUT_DATA = { 8'd0  ,2'b10,16'h3E54, 16'hEF00};
    391 : LUT_DATA = { 8'd0  ,2'b10,16'h3E55, 16'h1000};
    392 : LUT_DATA = { 8'd0  ,2'b10,16'h3E56, 16'hC000};
    393 : LUT_DATA = { 8'd0  ,2'b10,16'h3E57, 16'h6600};
    394 : LUT_DATA = { 8'd0  ,2'b10,16'h3E58, 16'h8500};
    395 : LUT_DATA = { 8'd0  ,2'b10,16'h3E59, 16'h6400};
    396 : LUT_DATA = { 8'd0  ,2'b10,16'h3E5A, 16'h8100};
    397 : LUT_DATA = { 8'd0  ,2'b10,16'h3E5B, 16'h1700};
    398 : LUT_DATA = { 8'd0  ,2'b10,16'h3E5C, 16'h0000};
    399 : LUT_DATA = { 8'd0  ,2'b10,16'h3E5D, 16'h8000};
    400 : LUT_DATA = { 8'd0  ,2'b10,16'h3E5E, 16'h2000};
    401 : LUT_DATA = { 8'd0  ,2'b10,16'h3E5F, 16'h0D00};
    402 : LUT_DATA = { 8'd0  ,2'b10,16'h3E60, 16'h8000};
    403 : LUT_DATA = { 8'd0  ,2'b10,16'h3E61, 16'h1800};
    404 : LUT_DATA = { 8'd0  ,2'b10,16'h3E62, 16'h0C00};
    405 : LUT_DATA = { 8'd0  ,2'b10,16'h3E63, 16'h8000};
    406 : LUT_DATA = { 8'd0  ,2'b10,16'h3E64, 16'h6400};
    407 : LUT_DATA = { 8'd0  ,2'b10,16'h3E65, 16'h3000};
    408 : LUT_DATA = { 8'd0  ,2'b10,16'h3E66, 16'h6000};
    409 : LUT_DATA = { 8'd0  ,2'b10,16'h3E67, 16'h4100};
    410 : LUT_DATA = { 8'd0  ,2'b10,16'h3E68, 16'h8200};
    411 : LUT_DATA = { 8'd0  ,2'b10,16'h3E69, 16'h4200};
    412 : LUT_DATA = { 8'd0  ,2'b10,16'h3E6A, 16'hB200};
    413 : LUT_DATA = { 8'd0  ,2'b10,16'h3E6B, 16'h4200};
    414 : LUT_DATA = { 8'd0  ,2'b10,16'h3E6C, 16'h8000};
    415 : LUT_DATA = { 8'd0  ,2'b10,16'h3E6D, 16'h4000};
    416 : LUT_DATA = { 8'd0  ,2'b10,16'h3E6E, 16'h8200};
    417 : LUT_DATA = { 8'd0  ,2'b10,16'h3E6F, 16'h4000};
    418 : LUT_DATA = { 8'd0  ,2'b10,16'h3E70, 16'h4C00};
    419 : LUT_DATA = { 8'd0  ,2'b10,16'h3E71, 16'h4500};
    420 : LUT_DATA = { 8'd0  ,2'b10,16'h3E72, 16'h9200};
    421 : LUT_DATA = { 8'd0  ,2'b10,16'h3E73, 16'h6A00};
    422 : LUT_DATA = { 8'd0  ,2'b10,16'h3E74, 16'h6B00};
    423 : LUT_DATA = { 8'd0  ,2'b10,16'h3E75, 16'h9B00};
    424 : LUT_DATA = { 8'd0  ,2'b10,16'h3E76, 16'h4500};
    425 : LUT_DATA = { 8'd0  ,2'b10,16'h3E77, 16'h8100};
    426 : LUT_DATA = { 8'd0  ,2'b10,16'h3E78, 16'h4C00};
    427 : LUT_DATA = { 8'd0  ,2'b10,16'h3E79, 16'h4000};
    428 : LUT_DATA = { 8'd0  ,2'b10,16'h3E7A, 16'h8C00};
    429 : LUT_DATA = { 8'd0  ,2'b10,16'h3E7B, 16'h3000};
    430 : LUT_DATA = { 8'd0  ,2'b10,16'h3E7C, 16'hA400};
    431 : LUT_DATA = { 8'd0  ,2'b10,16'h3E7D, 16'h6700};
    432 : LUT_DATA = { 8'd0  ,2'b10,16'h3E7E, 16'h8500};
    433 : LUT_DATA = { 8'd0  ,2'b10,16'h3E7F, 16'h6500};
    434 : LUT_DATA = { 8'd0  ,2'b10,16'h3E80, 16'h8700};
    435 : LUT_DATA = { 8'd0  ,2'b10,16'h3E81, 16'h6500};
    436 : LUT_DATA = { 8'd0  ,2'b10,16'h3E82, 16'h3000};
    437 : LUT_DATA = { 8'd0  ,2'b10,16'h3E83, 16'h6000};
    438 : LUT_DATA = { 8'd0  ,2'b10,16'h3E84, 16'hD300};
    439 : LUT_DATA = { 8'd0  ,2'b10,16'h3E85, 16'h6A00};
    440 : LUT_DATA = { 8'd0  ,2'b10,16'h3E86, 16'h6B00};
    441 : LUT_DATA = { 8'd0  ,2'b10,16'h3E87, 16'hAC00};
    442 : LUT_DATA = { 8'd0  ,2'b10,16'h3E88, 16'h6C00};
    443 : LUT_DATA = { 8'd0  ,2'b10,16'h3E89, 16'h3200};
    444 : LUT_DATA = { 8'd0  ,2'b10,16'h3E8A, 16'hA800};
    445 : LUT_DATA = { 8'd0  ,2'b10,16'h3E8B, 16'h8000};
    446 : LUT_DATA = { 8'd0  ,2'b10,16'h3E8C, 16'h2800};
    447 : LUT_DATA = { 8'd0  ,2'b10,16'h3E8D, 16'h3000};
    448 : LUT_DATA = { 8'd0  ,2'b10,16'h3E8E, 16'h7000};
    449 : LUT_DATA = { 8'd0  ,2'b10,16'h3E8F, 16'h0000};
    450 : LUT_DATA = { 8'd0  ,2'b10,16'h3E90, 16'h8000};
    451 : LUT_DATA = { 8'd0  ,2'b10,16'h3E91, 16'h4000};
    452 : LUT_DATA = { 8'd0  ,2'b10,16'h3E92, 16'h4C00};
    453 : LUT_DATA = { 8'd0  ,2'b10,16'h3E93, 16'hBD00};
    454 : LUT_DATA = { 8'd0  ,2'b10,16'h3E94, 16'h0000};
    455 : LUT_DATA = { 8'd0  ,2'b10,16'h3E95, 16'h0E00};
    456 : LUT_DATA = { 8'd0  ,2'b10,16'h3E96, 16'hBE00};
    457 : LUT_DATA = { 8'd0  ,2'b10,16'h3E97, 16'h4400};
    458 : LUT_DATA = { 8'd0  ,2'b10,16'h3E98, 16'h8800};
    459 : LUT_DATA = { 8'd0  ,2'b10,16'h3E99, 16'h4400};
    460 : LUT_DATA = { 8'd0  ,2'b10,16'h3E9A, 16'hBC00};
    461 : LUT_DATA = { 8'd0  ,2'b10,16'h3E9B, 16'h7800};
    462 : LUT_DATA = { 8'd0  ,2'b10,16'h3E9C, 16'h0900};
    463 : LUT_DATA = { 8'd0  ,2'b10,16'h3E9D, 16'h0000};
    464 : LUT_DATA = { 8'd0  ,2'b10,16'h3E9E, 16'h8900};
    465 : LUT_DATA = { 8'd0  ,2'b10,16'h3E9F, 16'h0400};
    466 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA0, 16'h8000};
    467 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA1, 16'h8000};
    468 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA2, 16'h0200};
    469 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA3, 16'h4000};
    470 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA4, 16'h8600};
    471 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA5, 16'h0900};
    472 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA6, 16'h0000};
    473 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA7, 16'h8E00};
    474 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA8, 16'h0900};
    475 : LUT_DATA = { 8'd0  ,2'b10,16'h3EA9, 16'h0000};
    476 : LUT_DATA = { 8'd0  ,2'b10,16'h3EAA, 16'h8000};
    477 : LUT_DATA = { 8'd0  ,2'b10,16'h3EAB, 16'h0200};
    478 : LUT_DATA = { 8'd0  ,2'b10,16'h3EAC, 16'h4000};
    479 : LUT_DATA = { 8'd0  ,2'b10,16'h3EAD, 16'h8000};
    480 : LUT_DATA = { 8'd0  ,2'b10,16'h3EAE, 16'h0400};
    481 : LUT_DATA = { 8'd0  ,2'b10,16'h3EAF, 16'h8000};
    482 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB0, 16'h8800};
    483 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB1, 16'h7D00};
    484 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB2, 16'h9E00};
    485 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB3, 16'h8600};
    486 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB4, 16'h0900};
    487 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB5, 16'h0000};
    488 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB6, 16'h8700};
    489 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB7, 16'h7A00};
    490 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB8, 16'h0000};
    491 : LUT_DATA = { 8'd0  ,2'b10,16'h3EB9, 16'h0E00};
    492 : LUT_DATA = { 8'd0  ,2'b10,16'h3EBA, 16'hC300};
    493 : LUT_DATA = { 8'd0  ,2'b10,16'h3EBB, 16'h7900};
    494 : LUT_DATA = { 8'd0  ,2'b10,16'h3EBC, 16'h4C00};
    495 : LUT_DATA = { 8'd0  ,2'b10,16'h3EBD, 16'h4000};
    496 : LUT_DATA = { 8'd0  ,2'b10,16'h3EBE, 16'hBF00};
    497 : LUT_DATA = { 8'd0  ,2'b10,16'h3EBF, 16'h7000};
    498 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC0, 16'h0000};
    499 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC1, 16'h0000};
    500 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC2, 16'h0000};
    501 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC3, 16'h0000};
    502 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC4, 16'h0000};
    503 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC5, 16'h0000};
    504 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC6, 16'h0000};
    505 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC7, 16'h0000};
    506 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC8, 16'h0000};
    507 : LUT_DATA = { 8'd0  ,2'b10,16'h3EC9, 16'h0000};
    508 : LUT_DATA = { 8'd0  ,2'b10,16'h3ECA, 16'h0000};
    509 : LUT_DATA = { 8'd0  ,2'b10,16'h3ECB, 16'h0000};
    510 : LUT_DATA = { 8'd0  ,2'b11,16'h301A, 16'h0018}; 	// RESET_REGISTER
    511 : LUT_DATA = { 8'd0  ,2'b11,16'h3EDE, 16'h6664}; 	// DAC_LD_18_19
    512 : LUT_DATA = { 8'd0  ,2'b11,16'h3EDE, 16'h6664}; 	// DAC_LD_18_19
    513 : LUT_DATA = { 8'd0  ,2'b11,16'h3EDE, 16'h6664}; 	// DAC_LD_18_19
    514 : LUT_DATA = { 8'd0  ,2'b11,16'h3EDE, 16'h6664}; 	// DAC_LD_18_19
    515 : LUT_DATA = { 8'd0  ,2'b11,16'h3EE0, 16'h26D5}; 	// DAC_LD_20_21
    516 : LUT_DATA = { 8'd0  ,2'b11,16'h3EE0, 16'h26D5}; 	// DAC_LD_20_21
    517 : LUT_DATA = { 8'd0  ,2'b11,16'h301A, 16'h001C}; 	// RESET_REGISTER
    518 : LUT_DATA = { 8'd0  ,2'b11,16'h0300, 16'h0005}; 	// VT_PIX_CLK_DIV
    519 : LUT_DATA = { 8'd0  ,2'b11,16'h0302, 16'h0001}; 	// VT_SYS_CLK_DIV
    520 : LUT_DATA = { 8'd0  ,2'b11,16'h0304, 16'h0004}; 	// PRE_PLL_CLK_DIV
    521 : LUT_DATA = { 8'd0  ,2'b11,16'h0306, 16'h007A}; 	// PLL_MULTIPLIER
    522 : LUT_DATA = { 8'd0  ,2'b11,16'h0308, 16'h000A}; 	// OP_PIX_CLK_DIV
    523 : LUT_DATA = { 8'd0  ,2'b11,16'h030A, 16'h0001}; 	// OP_SYS_CLK_DIV
    524 : LUT_DATA = { 8'd0  ,2'b11,16'h3064, 16'h7800}; 	// SMIA_TEST
    525 : LUT_DATA = { 8'd0  ,2'b11,16'h0300, 16'h0005}; 	// VT_PIX_CLK_DIV     // apply .ini from arrow, richard
    526 : LUT_DATA = { 8'd0  ,2'b11,16'h0302, 16'h0001}; 	// VT_SYS_CLK_DIV
    527 : LUT_DATA = { 8'd0  ,2'b11,16'h0304, 16'h0004}; 	// PRE_PLL_CLK_DIV
    528 : LUT_DATA = { 8'd0  ,2'b11,16'h0306, 16'h0046}; 	// PLL_MULTIPLIER
    529 : LUT_DATA = { 8'd0  ,2'b11,16'h0308, 16'h000A}; 	// OP_PIX_CLK_DIV
    530 : LUT_DATA = { 8'd0  ,2'b11,16'h030A, 16'h0001}; 	// OP_SYS_CLK_DIV     //VCO =  XTCLK * pll_multiplier(R0x306) / (pre_pll_clk_div(R0x0304)) = 24MHz * 0x46 / 4 = 24 * 70 / 4 = 420MHz// vt_sys_clk =  VCO / (vt_sys_clk_div(R0x302) x 2) = 420 / (1 x 2) = 210Mhz
    531 : LUT_DATA = { 8'd0  ,2'b11,16'h0300, 16'h0005}; 	// VT_PIX_CLK_DIV
    532 : LUT_DATA = { 8'd0  ,2'b11,16'h0302, 16'h0001}; 	// VT_SYS_CLK_DIV
    533 : LUT_DATA = { 8'd0  ,2'b11,16'h0304, 16'h0008}; 	// PRE_PLL_CLK_DIV
    534 : LUT_DATA = { 8'd0  ,2'b11,16'h0306, 16'h0046}; 	// PLL_MULTIPLIER
    535 : LUT_DATA = { 8'd0  ,2'b11,16'h0308, 16'h000A}; 	// OP_PIX_CLK_DIV
    536 : LUT_DATA = { 8'd0  ,2'b11,16'h030A, 16'h0001}; 	// OP_SYS_CLK_DIV    //VCO = 210MHz// vt_sys_clk = 105Mhz 
    537 : LUT_DATA = { 8'd0  ,2'b11,16'h0112, 16'h0808};        // CCP_DATA_FORMAT   // richard add: raw8
    538 : LUT_DATA = { 8'd1  ,2'b11,16'h31B0, 16'h0060}; 	// FRAME_PREAMBLE Sleep(1);
    539 : LUT_DATA = { 8'd0  ,2'b11,16'h31B2, 16'h0042}; 	// LINE_PREAMBLE
    540 : LUT_DATA = { 8'd0  ,2'b11,16'h31B4, 16'h1C36}; 	// MIPI_TIMING_0
    541 : LUT_DATA = { 8'd0  ,2'b11,16'h31B6, 16'h5218}; 	// MIPI_TIMING_1
    542 : LUT_DATA = { 8'd0  ,2'b11,16'h31B8, 16'h404A}; 	// MIPI_TIMING_2
    543 : LUT_DATA = { 8'd0  ,2'b11,16'h31BA, 16'h028A}; 	// MIPI_TIMING_3
    544 : LUT_DATA = { 8'd0  ,2'b11,16'h31BC, 16'h0008}; 	// MIPI_TIMING_4
    545 : LUT_DATA = { 8'd1  ,2'b11,16'h0342, 16'h1000}; 	// LINE_LENGTH_PCK  Sleep(1);
    546 : LUT_DATA = { 8'd0  ,2'b11,16'h0340, 16'h0556}; 	// FRAME_LENGTH_LINES
    547 : LUT_DATA = { 8'd0  ,2'b11,16'h0202, 16'h0500}; 	// COARSE_INTEGRATION_TIME
    548 : LUT_DATA = { 8'd0  ,2'b11,16'h0342, 16'h0ECE}; 	// LINE_LENGTH_PCK
    549 : LUT_DATA = { 8'd0  ,2'b11,16'h0340, 16'h0A0F}; 	// FRAME_LENGTH_LINES
    550 : LUT_DATA = { 8'd0  ,2'b11,16'h0202, 16'h0A0F}; 	// COARSE_INTEGRATION_TIME
   


    551 : LUT_DATA = {8'd0 ,2'b11, 16'h0344, 16'h0468}; 	// X_ADDR_START 0x0008+(3264-1024)/2 = 1128
    552 : LUT_DATA = {8'd0 ,2'b11, 16'h0348, 16'h0869}; 	// X_ADDR_END 8+1024+1+(3264-1024)/2 = 2153
    553 : LUT_DATA = {8'd0 ,2'b11, 16'h0346, 16'h0350}; 	// Y_ADDR_START 0x0008+(2448-768)/2 = 848
    554 : LUT_DATA = {8'd0 ,2'b11, 16'h034A, 16'h0651}; 	// Y_ADDR_END 8+768+1+(2448-768)/2 = 1617
	555 : LUT_DATA = {8'd0 ,2'b11, 16'h034C, 16'h0400}; 	// X_OUTPUT_SIZE
	556 : LUT_DATA = {8'd0 ,2'b11, 16'h034E, 16'h0300}; 	// Y_OUTPUT_SIZE
	557 : LUT_DATA = {8'd0 ,2'b11, 16'h020E, 16'h0100}; 	// digital_gain_greenr (default 0x100) // gain control (white balance)
	558 : LUT_DATA = {8'd0 ,2'b11, 16'h0210, 16'h0180}; 	// digital_gain_red (default 0x100)
	559 : LUT_DATA = {8'd0 ,2'b11, 16'h0212, 16'h0140}; 	// digital_gain_blue (default 0x100)
	560 : LUT_DATA = {8'd0 ,2'b11, 16'h0214, 16'h0100}; 	// digital_gain_greenb (default 0x100)
	561 : LUT_DATA = {8'd0 ,2'b11, 16'h3040, 16'h4041}; 	// READ_MODE
	562 : LUT_DATA = {8'd0 ,2'b11, 16'h3040, 16'h8041}; 	// READ_MODE
    563 : LUT_DATA = {8'd0 ,2'b11, 16'h0400, 16'h0000}; 	// SCALING_MODE, 0: disable scaling
	564 : LUT_DATA = {8'd0 ,2'b11, 16'h0402, 16'h0000}; 	// SPATIAL_SAMPLING
	565 : LUT_DATA = {8'd0 ,2'b11, 16'h0404, 16'h0020}; 	// SCALE_M (default 0x0010)
	566 : LUT_DATA = {8'd0 ,2'b11, 16'h0408, 16'h0208}; 	// SECOND_RESIDUAL
	567 : LUT_DATA = {8'd0 ,2'b11, 16'h040A, 16'h00C7}; 	// SECOND_CROP
	568 : LUT_DATA = {8'd0 ,2'b11, 16'h306E, 16'h9090}; 	// DATA_PATH_SELECT
	569 : LUT_DATA = {8'd0 ,2'b11, 16'h301A, 16'h001C}; 	// RESET_REGISTER (Lock_reg & stream)
//read	
	570 : LUT_DATA	=	{8'h0,2'b10,16'h0000, 16'h0};	//chip_version
	571 : LUT_DATA	=	{8'h0,2'b10,16'h0001, 16'h0};	
	572 : LUT_DATA	=	{8'h0,2'b10,16'h0002, 16'h0};   //revision_number
	573 : LUT_DATA	=	{8'h0,2'b10,16'h0003, 16'h0};   //manufacture_id
	574 : LUT_DATA	=	{8'h0,2'b10,16'h0004, 16'h0};   //smia_version
	      
	575 : LUT_DATA	=	{8'h10,2'b10,16'h0005,16'h0000};
	576 : LUT_DATA	=	{8'h10,2'b10,16'h0006,16'h0000};
	577 : LUT_DATA	=	{8'h10,2'b10,16'h0008,16'h0000};
	578 : LUT_DATA	=	{8'h10,2'b10,16'h0009,16'h0000};
	579 : LUT_DATA	=	{8'h10,2'b10,16'h3024,16'h0000};
	580 : LUT_DATA	=	{8'h10,2'b10,16'h3025,16'h0000};
	581 : LUT_DATA	=	{8'h10,2'b10,16'h0112,16'h0000};
	582 : LUT_DATA	=	{8'h10,2'b10,16'h0113,16'h0000};

	default:;
	endcase
end
endmodule
